lpm_compare1_inst : lpm_compare1 PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		AeB	 => AeB_sig,
		AlB	 => AlB_sig
	);
