lpm_dff1_inst : lpm_dff1 PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		q	 => q_sig
	);
