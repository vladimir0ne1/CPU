lpm_dff2_inst : lpm_dff2 PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		q	 => q_sig
	);
