lpm_counter1_inst : lpm_counter1 PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		sload	 => sload_sig,
		q	 => q_sig
	);
