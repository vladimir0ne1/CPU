lpm_compare4_inst : lpm_compare4 PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		AeB	 => AeB_sig,
		AgB	 => AgB_sig,
		AlB	 => AlB_sig
	);
