lpm_clshift0_inst : lpm_clshift0 PORT MAP (
		data	 => data_sig,
		distance	 => distance_sig,
		result	 => result_sig
	);
