lpm_bustri0_inst : lpm_bustri0 PORT MAP (
		data	 => data_sig,
		enabledt	 => enabledt_sig,
		tridata	 => tridata_sig
	);
