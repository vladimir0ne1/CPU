lpm_constant0_inst : lpm_constant0 PORT MAP (
		result	 => result_sig
	);
