lpm_compare3_inst : lpm_compare3 PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		AeB	 => AeB_sig
	);
