lpm_dff3_inst : lpm_dff3 PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		q	 => q_sig
	);
