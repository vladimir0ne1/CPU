lpm_dff0_inst : lpm_dff0 PORT MAP (
		clock	 => clock_sig,
		data	 => data_sig,
		q	 => q_sig
	);
